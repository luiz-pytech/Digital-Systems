entity Cambio_Automatico is
port(
  s : in bit

);

end Cambio_Automatico;

architecture behav of Cambio_Automatico is
begin


end architecture behav;